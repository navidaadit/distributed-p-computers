`timescale 1ns / 1ps
module LUT_bias ( Iin, Out);

import PSL_pkg :: *;

input  [i_bit_width-2:0] Iin;
output reg [RNG_bit_width-1:0] Out;

always @ *//( posedge En )
begin 
case (Iin)

5'b00000 : Out =32'b10000000000000000000000000000000;
5'b00001 : Out =32'b10111011001001101010011110101111;
5'b00010 : Out =32'b11100001011110111110101011010100;
5'b00011 : Out =32'b11110011110110111110010111100010;
5'b00100 : Out =32'b11111011011001010100000101111000;
5'b00101 : Out =32'b11111110010010010110000010011000;
5'b00110 : Out =32'b11111111010111011111010001000100;
5'b00111 : Out =32'b11111111110001000100101100011001;
5'b01000 : Out =32'b11111111111010100000010111000010;
5'b01001 : Out =32'b11111111111101111110100111001000;
5'b01010 : Out =32'b11111111111111010000011001011010;
5'b01011 : Out =32'b11111111111111101110011111001100;
5'b01100 : Out =32'b11111111111111111001100011101011;
5'b01101 : Out =32'b11111111111111111101101000010100;
5'b01110 : Out =32'b11111111111111111111001000001101;
5'b01111 : Out =32'b11111111111111111111101011011110;
5'b10000 : Out =32'b11111111111111111111111000011101;
5'b10001 : Out =32'b11111111111111111111111101001110;
5'b10010 : Out =32'b11111111111111111111111110111111;
5'b10011 : Out =32'b11111111111111111111111111101000;
5'b10100 : Out =32'b11111111111111111111111111110111;
5'b10101 : Out =32'b11111111111111111111111111111101;
5'b10110 : Out =32'b11111111111111111111111111111111;
5'b10111 : Out =32'b11111111111111111111111111111111;
5'b11000 : Out =32'b11111111111111111111111111111111;
5'b11001 : Out =32'b11111111111111111111111111111111;
5'b11010 : Out =32'b11111111111111111111111111111111;
5'b11011 : Out =32'b11111111111111111111111111111111;
5'b11100 : Out =32'b11111111111111111111111111111111;
5'b11101 : Out =32'b11111111111111111111111111111111;
5'b11110 : Out =32'b11111111111111111111111111111111;
5'b11111 : Out =32'b11111111111111111111111111111111;

endcase
end
endmodule